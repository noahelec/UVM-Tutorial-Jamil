interface our_interface(input logic clk);
    //input_1
    //input_2

    //output

    logic [7:0] input_1;
    logic [7:0] input_2;

    logic [15:0] output_3;
endinterface //